`timescale 1ns / 1ps

`include "global.vh"

module CPU_tb;

logic CLK,UART_RX,INITIALIZE,START_EXEC,UART_TX;
logic[7:0] LED;
CPU CPU(.*);

parameter INST_LEN = 318;
logic[31:0] data[INST_LEN] = {
32'b00000000000000000000000000000000,
32'b10111111100000000000000000000000,
32'b10111111110000000000000000000000,
32'b00111110010011001100110011001101,
32'b01000000100000000000000000000000,
32'b11001011000000000000000000000000,
32'b01001011000000000000000000000000,
32'b00000000011111111111111111111111,
32'b01001011000000000000000000000000,
32'b00000000100000000000000000000000,
32'b00000000100000000000000000000000,
32'b00000000100000000000000000000000,
32'b11111111111111111111111111111111,
32'b01001111100001001110001000000000, // Li (Reg 28) (Imm 10000)
32'b01001100000000000000000000000000, // Li (Reg 0) (Imm 0)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01001100010000000000101000000000, // Li (Reg 2) (Imm 80)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000011000100000, // Li (Reg 2) (Imm 49)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000000101000000, // Li (Reg 2) (Imm 10)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000011010100000, // Li (Reg 2) (Imm 53)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000010000000000, // Li (Reg 2) (Imm 32)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000011010100000, // Li (Reg 2) (Imm 53)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000000101000000, // Li (Reg 2) (Imm 10)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b01001100010000000000000000000000, // Li (Reg 2) (Imm 0)
32'b11111100010001000000000000110111, // Bgti (Reg 2) (Imm5 4) (LabelI "yloop.604.exit.1075")
32'b01001100011000000000000000000000, // Li (Reg 3) (Imm 0)
32'b01100100010111010000000000000001, // Sw (Reg 2) (Reg 29) (Imm 1)
32'b11001100010000110000000000000000, // Swap (Reg 2) (Reg 3)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000101101010000000000, // Jal (LabelI "xloop.607")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b01011000010111010000000000000001, // Lwr (Reg 2) (Reg 29) (Imm 1)
32'b00010000010000100000000000000001, // Addi (Reg 2) (Reg 2) (Imm 1)
32'b10001000000000001011010000000000, // J (LabelI "tailrecurse.i.1075")
32'b11001000000000000000000000000000, // Exit
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11110100010000010000000000111100, // Bnei (Reg 2) (Imm5 1) (LabelI "else.989.1084")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01011100001000000000000011000000, // Lsl (FReg 1) (LabelF "l.1086")
32'b00110100000000010000000000000000, // Adds (FReg 0) (FReg 1) (FReg 0)
32'b00010000010000101111111111111111, // Addi (Reg 2) (Reg 2) (Imm (-1))
32'b10001000000000001110010000000000, // J (LabelI "tailrecurse.1084")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01111000010000110000000001000100, // Bgt (Reg 2) (Reg 3) (LabelI "else.994.1087")
32'b10011100010000100000000000000001, // Slli (Reg 2) (Reg 2) (Imm 1)
32'b10001000000000010000010000000000, // J (LabelI "tailrecurse.1087")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01111000011001000000000001001111, // Bgt (Reg 3) (Reg 4) (LabelI "else.999.1088")
32'b00101000101000100000000000000010, // Divi (Reg 5) (Reg 2) (Imm 2)
32'b01110100100000100000000001001101, // Blt (Reg 4) (Reg 2) (LabelI "else.1002.1088")
32'b00010100100001000001000000000000, // Sub (Reg 4) (Reg 4) (Reg 2)
32'b00000100010001010000000000000000, // Move (Reg 2) (Reg 5)
32'b10001000000000010001110000000000, // J (LabelI "tailrecurse.1088")
32'b00000100010001010000000000000000, // Move (Reg 2) (Reg 5)
32'b10001000000000010001110000000000, // J (LabelI "tailrecurse.1088")
32'b00000100010001000000000000000000, // Move (Reg 2) (Reg 4)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11100000101000101111110100000000, // Cmpi GT (Reg 5) (Reg 2) (Imm5 (-1))
32'b00001000011000100000000000000000, // Neg (Reg 3) (Reg 2)
32'b11010100011001010001000011000000, // Select (Reg 3) (Reg 5) (Reg 2) (Reg 3)
32'b01010111011000000000000011100000, // Lwl (Reg 27) (LabelF "bigint.7")
32'b01111000011110110000000001100101, // Bgt (Reg 3) (Reg 27) (LabelI "then.1013.1089")
32'b01010111011000000000000100000000, // Lwl (Reg 27) (LabelF "bigint.8")
32'b00001100010000111101100000000000, // Add (Reg 2) (Reg 3) (Reg 27)
32'b11101000000000100000000000000000, // Cvtsw (FReg 0) (Reg 2)
32'b01011100001000000000000010100000, // Lsl (FReg 1) (LabelF "l.1093")
32'b00110100000000010000000000000000, // Adds (FReg 0) (FReg 1) (FReg 0)
32'b10101100101000010000000001011111, // Beqi (Reg 5) (Imm5 1) (LabelI "phi_else.1014.1089_then.1016.1089")
32'b10001000000000011000010000000000, // J (LabelI "else.1021.1089")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b00110000001000000000000000000000, // Negs (FReg 1) (FReg 0)
32'b00101100000000010000000000000000, // Movs (FReg 0) (FReg 1)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01010111011000000000000100100000, // Lwl (Reg 27) (LabelF "bigint.9")
32'b00100100010000111101100000000000, // Div (Reg 2) (Reg 3) (Reg 27)
32'b01010111011000000000000101000000, // Lwl (Reg 27) (LabelF "bigint.10")
32'b00000100100110110000000000000000, // Move (Reg 4) (Reg 27)
32'b01111000100000110000000001101100, // Bgt (Reg 4) (Reg 3) (LabelI "sub1_mod.536.exit.1089")
32'b10011100100001000000000000000001, // Slli (Reg 4) (Reg 4) (Imm 1)
32'b10001000000000011010010000000000, // J (LabelI "tailrecurse.i.1089")
32'b01010111011000000000000101100000, // Lwl (Reg 27) (LabelF "bigint.11")
32'b00000100110110110000000000000000, // Move (Reg 6) (Reg 27)
32'b01111000110000110000000001110110, // Bgt (Reg 6) (Reg 3) (LabelI "sub2_mod.541.exit.1089")
32'b00101000110001000000000000000010, // Divi (Reg 6) (Reg 4) (Imm 2)
32'b01110100011001000000000001110100, // Blt (Reg 3) (Reg 4) (LabelI "else.1002.i.1089")
32'b00010100011000110010000000000000, // Sub (Reg 3) (Reg 3) (Reg 4)
32'b00000100100001100000000000000000, // Move (Reg 4) (Reg 6)
32'b10001000000000011011000000000000, // J (LabelI "tailrecurse.i1.1089")
32'b00000100100001100000000000000000, // Move (Reg 4) (Reg 6)
32'b10001000000000011011000000000000, // J (LabelI "tailrecurse.i1.1089")
32'b01011100000000000000000011000000, // Lsl (FReg 0) (LabelF "l.1086")
32'b11110100010000010000000010001000, // Bnei (Reg 2) (Imm5 1) (LabelI "else.989.i.1089")
32'b01100100101111010000000000000001, // Sw (Reg 5) (Reg 29) (Imm 1)
32'b01101000000111010000000000000010, // Ss (FReg 0) (Reg 29) (Imm 2)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000011, // Addi (Reg 29) (Reg 29) (Imm 3)
32'b10010000000000010100100000000000, // Jal (LabelI "float_of_int.554")
32'b00010011101111011111111111111101, // Addi (Reg 29) (Reg 29) (Imm (-3))
32'b00101100001000000000000000000000, // Movs (FReg 1) (FReg 0)
32'b01100000000111010000000000000010, // Lsr (FReg 0) (Reg 29) (Imm 2)
32'b00110100000000000000100000000000, // Adds (FReg 0) (FReg 0) (FReg 1)
32'b01011000101111010000000000000001, // Lwr (Reg 5) (Reg 29) (Imm 1)
32'b10101100101000010000000010000100, // Beqi (Reg 5) (Imm5 1) (LabelI "phi_iaf_mul.490.exit.1089_then.1016.1089")
32'b10001000000000100001010000000000, // J (LabelI "else.1017.1089")
32'b10001000000000010111110000000000, // J (LabelI "then.1016.1089")
32'b00110000000000000000000000000000, // Negs (FReg 0) (FReg 0)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01011100001000000000000011000000, // Lsl (FReg 1) (LabelF "l.1086")
32'b00110100000000010000000000000000, // Adds (FReg 0) (FReg 1) (FReg 0)
32'b00010000010000101111111111111111, // Addi (Reg 2) (Reg 2) (Imm (-1))
32'b10001000000000011101110000000000, // J (LabelI "tailrecurse.i2.1089")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11111100010010010000000010010001, // Bgti (Reg 2) (Imm5 9) (LabelI "then.1025.1094")
32'b00010000010000100000000000110000, // Addi (Reg 2) (Reg 2) (Imm 48)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000001000101000000000000, // J (LabelI "min_caml_print_char")
32'b00101000011000100000000000001010, // Divi (Reg 3) (Reg 2) (Imm 10)
32'b01100100011111010000000000000001, // Sw (Reg 3) (Reg 29) (Imm 1)
32'b01100100010111010000000000000010, // Sw (Reg 2) (Reg 29) (Imm 2)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000011, // Addi (Reg 29) (Reg 29) (Imm 3)
32'b10010000000000100011000000000000, // Jal (LabelI "print_int_sub.296.887")
32'b00010011101111011111111111111101, // Addi (Reg 29) (Reg 29) (Imm (-3))
32'b01011000011111010000000000000001, // Lwr (Reg 3) (Reg 29) (Imm 1)
32'b00100000011000111111111111110110, // Multi (Reg 3) (Reg 3) (Imm (-10))
32'b01011000010111010000000000000010, // Lwr (Reg 2) (Reg 29) (Imm 2)
32'b00010000010000100000000000110000, // Addi (Reg 2) (Reg 2) (Imm 48)
32'b00001100010000100001100000000000, // Add (Reg 2) (Reg 2) (Reg 3)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000001000101000000000000, // J (LabelI "min_caml_print_char")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11010000000000100000000000000000, // Swaps (FReg 0) (FReg 2)
32'b11110100010000000000000010100101, // Bnei (Reg 2) (Imm5 0) (LabelI "else.1056.1095")
32'b01001100010000000000011000100000, // Li (Reg 2) (Imm 49)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000001000101000000000000, // J (LabelI "min_caml_print_char")
32'b00111000011000000001100000000000, // Subs (FReg 3) (FReg 0) (FReg 3)
32'b00110100011000110010000000000000, // Adds (FReg 3) (FReg 3) (FReg 4)
32'b00110100010000100001000000000000, // Adds (FReg 2) (FReg 2) (FReg 2)
32'b00111100010000100000100000000000, // Muls (FReg 2) (FReg 2) (FReg 1)
32'b00110100001000100010100000000000, // Adds (FReg 1) (FReg 2) (FReg 5)
32'b00111100000000110001100000000000, // Muls (FReg 0) (FReg 3) (FReg 3)
32'b00111100010000010000100000000000, // Muls (FReg 2) (FReg 1) (FReg 1)
32'b00110100110000000001000000000000, // Adds (FReg 6) (FReg 0) (FReg 2)
32'b01011100111000000000000010000000, // Lsl (FReg 7) (LabelF "l.1098")
32'b10000000110001110000000010110010, // Cles (FReg 6) (FReg 7) (LabelI "then.1059.1095")
32'b01001100010000000000011000000000, // Li (Reg 2) (Imm 48)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000001000101000000000000, // J (LabelI "min_caml_print_char")
32'b00010000010000101111111111111111, // Addi (Reg 2) (Reg 2) (Imm (-1))
32'b11010000011000100000000000000000, // Swaps (FReg 3) (FReg 2)
32'b10001000000000101000010000000000, // J (LabelI "tailrecurse.1095")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b11111100100001000000000011111001, // Bgti (Reg 4) (Imm5 4) (LabelI "then.1065.1100")
32'b01100100100111010000000000000001, // Sw (Reg 4) (Reg 29) (Imm 1)
32'b01100100011111010000000000000010, // Sw (Reg 3) (Reg 29) (Imm 2)
32'b00000100010001000000000000000000, // Move (Reg 2) (Reg 4)
32'b00010011101111010000000000000011, // Addi (Reg 29) (Reg 29) (Imm 3)
32'b10010000000000010100100000000000, // Jal (LabelI "float_of_int.554")
32'b00010011101111011111111111111101, // Addi (Reg 29) (Reg 29) (Imm (-3))
32'b00110100000000000000000000000000, // Adds (FReg 0) (FReg 0) (FReg 0)
32'b01011100001000000000000001100000, // Lsl (FReg 1) (LabelF "l.1102")
32'b00111100001000010000000000000000, // Muls (FReg 1) (FReg 1) (FReg 0)
32'b01011100000000000000000001000000, // Lsl (FReg 0) (LabelF "l.1104")
32'b00110100010000000000100000000000, // Adds (FReg 2) (FReg 0) (FReg 1)
32'b01101000010111010000000000000011, // Ss (FReg 2) (Reg 29) (Imm 3)
32'b01011000011111010000000000000010, // Lwr (Reg 3) (Reg 29) (Imm 2)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000100, // Addi (Reg 29) (Reg 29) (Imm 4)
32'b10010000000000010100100000000000, // Jal (LabelI "float_of_int.554")
32'b00010011101111011111111111111100, // Addi (Reg 29) (Reg 29) (Imm (-4))
32'b00101100001000000000000000000000, // Movs (FReg 1) (FReg 0)
32'b00110100001000010000100000000000, // Adds (FReg 1) (FReg 1) (FReg 1)
32'b01011100000000000000000001100000, // Lsl (FReg 0) (LabelF "l.1102")
32'b00111100000000000000100000000000, // Muls (FReg 0) (FReg 0) (FReg 1)
32'b01011100001000000000000000100000, // Lsl (FReg 1) (LabelF "l.1107")
32'b00110100001000010000000000000000, // Adds (FReg 1) (FReg 1) (FReg 0)
32'b01011000100111010000000000000001, // Lwr (Reg 4) (Reg 29) (Imm 1)
32'b01011000011111010000000000000010, // Lwr (Reg 3) (Reg 29) (Imm 2)
32'b01100000010111010000000000000011, // Lsr (FReg 2) (Reg 29) (Imm 3)
32'b01001100010000000000000000100000, // Li (Reg 2) (Imm 1)
32'b01011100110000000000000000000000, // Lsl (FReg 6) (LabelF "l.1108")
32'b01011100011000000000000000000000, // Lsl (FReg 3) (LabelF "l.1108")
32'b01011100000000000000000000000000, // Lsl (FReg 0) (LabelF "l.1108")
32'b01011100100000000000000000000000, // Lsl (FReg 4) (LabelF "l.1108")
32'b11110100010000000000000011100011, // Bnei (Reg 2) (Imm5 0) (LabelI "else.1056.i.1100")
32'b01001100010000000000011000100000, // Li (Reg 2) (Imm 49)
32'b01100100100111010000000000000001, // Sw (Reg 4) (Reg 29) (Imm 1)
32'b01100100011111010000000000000010, // Sw (Reg 3) (Reg 29) (Imm 2)
32'b00010011101111010000000000000100, // Addi (Reg 29) (Reg 29) (Imm 4)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111100, // Addi (Reg 29) (Reg 29) (Imm (-4))
32'b01011000100111010000000000000001, // Lwr (Reg 4) (Reg 29) (Imm 1)
32'b01011000011111010000000000000010, // Lwr (Reg 3) (Reg 29) (Imm 2)
32'b00010000010001000000000000000001, // Addi (Reg 2) (Reg 4) (Imm 1)
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b10001000000000101101110000000000, // J (LabelI "tailrecurse.1100")
32'b00111000101000110011000000000000, // Subs (FReg 5) (FReg 3) (FReg 6)
32'b00110100101001010001000000000000, // Adds (FReg 5) (FReg 5) (FReg 2)
32'b00110100100001000010000000000000, // Adds (FReg 4) (FReg 4) (FReg 4)
32'b00111100000001000000000000000000, // Muls (FReg 0) (FReg 4) (FReg 0)
32'b00110100000000000000100000000000, // Adds (FReg 0) (FReg 0) (FReg 1)
32'b00111100011001010010100000000000, // Muls (FReg 3) (FReg 5) (FReg 5)
32'b00111100110000000000000000000000, // Muls (FReg 6) (FReg 0) (FReg 0)
32'b00110100100000110011000000000000, // Adds (FReg 4) (FReg 3) (FReg 6)
32'b01011100111000000000000010000000, // Lsl (FReg 7) (LabelF "l.1098")
32'b10000000100001110000000011110110, // Cles (FReg 4) (FReg 7) (LabelI "then.1059.i.1100")
32'b01001100010000000000011000000000, // Li (Reg 2) (Imm 48)
32'b01100100100111010000000000000001, // Sw (Reg 4) (Reg 29) (Imm 1)
32'b01100100011111010000000000000010, // Sw (Reg 3) (Reg 29) (Imm 2)
32'b00010011101111010000000000000100, // Addi (Reg 29) (Reg 29) (Imm 4)
32'b10010000000001000101000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111100, // Addi (Reg 29) (Reg 29) (Imm (-4))
32'b01011000100111010000000000000001, // Lwr (Reg 4) (Reg 29) (Imm 1)
32'b01011000011111010000000000000010, // Lwr (Reg 3) (Reg 29) (Imm 2)
32'b10001000000000111000000000000000, // J (LabelI "iloop.623.exit.1100")
32'b00010000010000101111111111111111, // Addi (Reg 2) (Reg 2) (Imm (-1))
32'b00101100100001010000000000000000, // Movs (FReg 4) (FReg 5)
32'b10001000000000110101110000000000, // J (LabelI "tailrecurse.i.1100")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11111100010001000000000100000110, // Bgti (Reg 2) (Imm5 4) (LabelI "then.1070.1112")
32'b01001100011000000000000000000000, // Li (Reg 3) (Imm 0)
32'b01100100010111010000000000000001, // Sw (Reg 2) (Reg 29) (Imm 1)
32'b11001100010000110000000000000000, // Swap (Reg 2) (Reg 3)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000101101010000000000, // Jal (LabelI "xloop.607")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b01011000010111010000000000000001, // Lwr (Reg 2) (Reg 29) (Imm 1)
32'b00010000010000100000000000000001, // Addi (Reg 2) (Reg 2) (Imm 1)
32'b10001000000000111111000000000000, // J (LabelI "tailrecurse.1112")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000100011000000000000, // J (LabelI "print_int_sub.296.887")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000100011000000000000, // J (LabelI "print_int_sub.296.887")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000100011000000000000, // J (LabelI "print_int_sub.296.887")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000100011000000000000, // J (LabelI "print_int_sub.296.887")
32'b10100000010000000000000000000000, // PrintC (Reg 2)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b10100100010000000000000000000000, // ReadI (Reg 2)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b10101000000000000000000000000000, // ReadF (FReg 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b00000100110000100000000000000000, // Move (Reg 6) (Reg 2)
32'b01001100101000000000000000000000, // Li (Reg 5) (Imm 0)
32'b01110000011001010000000100011110, // Bne (Reg 3) (Reg 5) (LabelI "min_caml_init_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100100100001100000000000000000, // Sw (Reg 4) (Reg 6) (Imm 0)
32'b00010000011000111111111111111111, // Addi (Reg 3) (Reg 3) (Imm (-1))
32'b00010000110001100000000000000001, // Addi (Reg 6) (Reg 6) (Imm 1)
32'b10001000000001000111000000000000, // J (LabelI "min_caml_init_array_loop")
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b00000100010111000000000000000000, // Move (Reg 2) (Reg 28)
32'b01001100110000000000000000000000, // Li (Reg 6) (Imm 0)
32'b01110000100001100000000100100111, // Bne (Reg 4) (Reg 6) (LabelI "min_caml_create_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100100011111000000000000000000, // Sw (Reg 3) (Reg 28) (Imm 0)
32'b00010000100001001111111111111111, // Addi (Reg 4) (Reg 4) (Imm (-1))
32'b00010011100111000000000000000001, // Addi (Reg 28) (Reg 28) (Imm 1)
32'b10001000000001001001010000000000, // J (LabelI "min_caml_create_array_loop")
32'b00000100110000100000000000000000, // Move (Reg 6) (Reg 2)
32'b01001100101000000000000000000000, // Li (Reg 5) (Imm 0)
32'b01110000011001010000000100101111, // Bne (Reg 3) (Reg 5) (LabelI "min_caml_init_float_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01101000000001100000000000000000, // Ss (FReg 0) (Reg 6) (Imm 0)
32'b00010000011000111111111111111111, // Addi (Reg 3) (Reg 3) (Imm (-1))
32'b00010000110001100000000000000001, // Addi (Reg 6) (Reg 6) (Imm 1)
32'b10001000000001001011010000000000, // J (LabelI "min_caml_init_float_array_loop")
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b00000100010111000000000000000000, // Move (Reg 2) (Reg 28)
32'b01001100110000000000000000000000, // Li (Reg 6) (Imm 0)
32'b01110000100001100000000100111000, // Bne (Reg 4) (Reg 6) (LabelI "min_caml_create_float_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01101000000111000000000000000000, // Ss (FReg 0) (Reg 28) (Imm 0)
32'b00010000100001001111111111111111, // Addi (Reg 4) (Reg 4) (Imm (-1))
32'b00010011100111000000000000000001, // Addi (Reg 28) (Reg 28) (Imm 1)
32'b10001000000001001101100000000000, // J (LabelI "min_caml_create_float_array_loop")
32'b00000000000000000000000000000000, // Sqrt (FReg 0) (FReg 0)
32'b10001111111000000000000000000000 // Jr (Reg 31)
};
logic[9:0] in;
integer inst_itr;
integer byte_itr;
integer bit_itr;

initial begin
	CLK = 0;
	inst_itr = 0;
	byte_itr = 0;
	INITIALIZE <= 1;
	@(posedge CLK);
	INITIALIZE <= 0;
	repeat(INST_LEN) begin
		byte_itr = 0;
		repeat(4) begin
			unique case (byte_itr)
				0: in = {1'b1,data[inst_itr][31:24],1'b0};
				1: in = {1'b1,data[inst_itr][23:16],1'b0};
				2: in = {1'b1,data[inst_itr][15:8],1'b0};
				3: in = {1'b1,data[inst_itr][7:0],1'b0};
			endcase
			bit_itr = 0;
			repeat(10) begin
				UART_RX = in[bit_itr];
				repeat(T) @(posedge CLK);
				bit_itr = bit_itr + 1;
			end
			byte_itr = byte_itr + 1;
		end
		inst_itr = inst_itr + 1;
	end
	repeat(100) @(posedge CLK);
	START_EXEC = 1;
	repeat(2) @(posedge CLK);
	START_EXEC = 0;
end

always begin
	#33.3ns CLK=~CLK;
end

endmodule