`timescale 1ns / 1ps

parameter T=2604;

module CPU_tb;

logic CLK,UART_RX,INITIALIZE,START_EXEC,UART_TX;
logic[0:0] LED;
CPU CPU(.*);

parameter INST_LEN = 146;
logic[31:0] data[INST_LEN] = {
//32'b01010011110100110101001111110111,		//float
//32'b11111111111111111111111111111111,		//delimiter
//32'b010011_00000_0000000000000000_11010,	//li 0 0
//32'b000100_00000_00000_1000000000000010,	//addi 0 0 -hoge
//32'b010011_00001_1000000000000001_11010,	//li 1 10..01
//32'b000001_00010_00001_0101001101010111, 	//mv to 2 from 1
//32'b000010_00010_00001_0101001101010111, 	//neg 2 1
//32'b100110_00010_000010101001101010111, 	//print reg[2]
//32'b110010_00010000010101001101010111 	//exit
32'b00000000000000000000000000000000,
32'b10000000000000000000000000000000,
32'b00111111100000000000000000000000,
32'b01000000000000000000000000000000,
32'b00111111000000000000000000000000,
32'b01000000010010010000111111011011,
32'b00111111110010010000111111011011,
32'b11111111111111111111111111111111,
32'b01100111111111010000000000000001,
32'b01100111110111010000000000000010,
32'b00010011101111010000000000000110,
32'b00010011110111010000000000000000,
32'b01001100010000000000001010000000,
32'b01100111111111010000000000000000,
32'b00010011101111010000000000000001,
32'b10010000000000000101010000000000,
32'b00010011101111011111111111111111,
32'b01011011111111010000000000000000,
32'b01100111111111010000000000000000,
32'b00010011101111010000000000000001,
32'b10010000000000001011110000000000,
32'b00010011101111011111111111111111,
32'b01011011111111010000000000000000,
32'b00000111101111100000000000000000,
32'b00011011101111010000000000000110,
32'b01011011111111010000000000000001,
32'b01011011110111010000000000000010,
32'b01001100010000000000000000000000,
32'b11001000000000000000000000000000,
32'b01001100011000000000000000100000,
32'b01111000010000110000000000011000,
32'b10001111111000000000000000000000,
32'b00010000011000101111111111111111,
32'b01100100010111010000000000000000,
32'b00010000010000110000000000000000,
32'b01100111111111010000000000000001,
32'b00010011101111010000000000000010,
32'b10010000000000000101010000000000,
32'b00010011101111011111111111111110,
32'b01011011111111010000000000000001,
32'b01011000011111010000000000000000,
32'b00010000011000111111111111111110,
32'b01100100010111010000000000000001,
32'b00010000010000110000000000000000,
32'b01100111111111010000000000000010,
32'b00010011101111010000000000000011,
32'b10010000000000000101010000000000,
32'b00010011101111011111111111111101,
32'b01011011111111010000000000000010,
32'b01011000011111010000000000000001,
32'b00001100010000110001000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000101000000,
32'b10100000010000000000000000000000,
32'b10001111111000000000000000000000,
32'b10011000010000000000000000000000,
32'b10001111111000000000000000000000,
32'b10100000010000000000000000000000,
32'b10001111111000000000000000000000,
32'b10011100000000000000000000000000,
32'b10001111111000000000000000000000,
32'b10100100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b10101000000000000000000000000000,
32'b10001111111000000000000000000000,
32'b00000100100000100000000000000000,
32'b00000100010111000000000000000000,
32'b01001100110000000000000000000000,
32'b01110000100001100000000000111110,
32'b10001111111000000000000000000000,
32'b01100100011111000000000000000000,
32'b00010000100001001111111111111111,
32'b00010011100111000000000000000100,
32'b10001000000000001110110000000000,
32'b00000100100000100000000000000000,
32'b00000100010111000000000000000000,
32'b01001100110000000000000000000000,
32'b01110000100001100000000001000111,
32'b10001111111000000000000000000000,
32'b01101000000111000000000000000000,
32'b00010000100001001111111111111111,
32'b00010011100111000000000000000100,
32'b10001000000000010001000000000000,
32'b10001000000000010011000000000000,
32'b11000000010000000000000000000000,
32'b10001111111000000000000000000000,
32'b11000100000000100000000000000000,
32'b10001111111000000000000000000000,
32'b10111000000000000000000000000000,
32'b10001111111000000000000000000000,
32'b10111100000000000000000000000000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000000000000,
32'b01111100000000010000000001011010,
32'b01011100001000000000000000100000,
32'b01111100000000010000000001011010,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000000000000,
32'b10000100001000000000000001100000,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000000000000,
32'b10000100000000010000000001100000,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01001100100000000000000000000000,
32'b01101100010001000000000001101111,
32'b01101100011001000000000001101101,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01101100011001000000000001110010,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b10000100000000010000000001110111,
32'b01001100010000000000000000000000,
32'b10001111111000000000000000000000,
32'b01001100010000000000000000100000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000000000000,
32'b00111000000000010000000000000000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000000000000,
32'b10000100000000010000000001111001,
32'b10001111111000000000000000000000,
32'b00111100000000000000000000000000,
32'b10001111111000000000000000000000,
32'b01011100001000000000000010000000,
32'b00111100000000000000100000000000,
32'b10001111111000000000000000000000,
32'b10101100000000000000000000000000,
32'b10001111111000000000000000000000,
32'b10110000000000000000000000000000,
32'b10001111111000000000000000000000,
32'b10110100000000000000000000000000,
32'b10001111111000000000000000000000
};
logic[9:0] in;
integer inst_itr;
integer byte_itr;
integer bit_itr;

initial begin
	CLK = 0;
	inst_itr = 0;
	byte_itr = 0;
	INITIALIZE <= 1;
	@(posedge CLK);
	INITIALIZE <= 0;
	repeat(INST_LEN) begin
		byte_itr = 0;
		repeat(4) begin
			unique case (byte_itr)
				0: in = {1'b1,data[inst_itr][31:24],1'b0};
				1: in = {1'b1,data[inst_itr][23:16],1'b0};
				2: in = {1'b1,data[inst_itr][15:8],1'b0};
				3: in = {1'b1,data[inst_itr][7:0],1'b0};
			endcase
			bit_itr = 0;
			repeat(10) begin
				UART_RX = in[bit_itr];
				repeat(T) @(posedge CLK);
				bit_itr = bit_itr + 1;
			end
			byte_itr = byte_itr + 1;
		end
		inst_itr = inst_itr + 1;
	end
	repeat(100) @(posedge CLK);
	START_EXEC = 1;
	repeat(2) @(posedge CLK);
	START_EXEC = 0;
end

always begin
	#1ns CLK=~CLK;
end

endmodule