`define global
