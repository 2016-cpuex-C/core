`timescale 1ns / 1ps

`include "global.vh"

module CPU_tb;

logic CLK,UART_RX,INITIALIZE,START_EXEC,UART_TX;
logic[7:0] LED;
CPU CPU(.*);

parameter INST_LEN = 122;
logic[31:0] data[INST_LEN] = {
32'b11111111111111111111111111111111,
32'b01001111100001001110001000000000, // Li (Reg 28) (Imm 10000)
32'b01001100000000000000000000000000, // Li (Reg 0) (Imm 0)
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b01001100010000000000000010000000, // Li (Reg 2) (Imm 4)
32'b00010011101111010000000000000001, // Addi (Reg 29) (Reg 29) (Imm 1)
32'b10010000000000001110100000000000, // Jal (LabelI "fib.707")
32'b00010011101111011111111111111111, // Addi (Reg 29) (Reg 29) (Imm (-1))
32'b11111100010111110000000000010101, // Bgti (Reg 2) (Imm5 (-1)) (LabelI "then.728.i.738")
32'b01001100011000000000010110100000, // Li (Reg 3) (Imm 45)
32'b01100100010111010000000000000001, // Sw (Reg 2) (Reg 29) (Imm 1)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000010100000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b01011000010111010000000000000001, // Lwr (Reg 2) (Reg 29) (Imm 1)
32'b00001000010000100000000000000000, // Neg (Reg 2) (Reg 2)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000000110010000000000, // Jal (LabelI "print_int_sub.328")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b11001000000000000000000000000000, // Exit
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000000110010000000000, // Jal (LabelI "print_int_sub.328")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b10001000000000000101000000000000, // J (LabelI "print_int.326.exit.738")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11111100010010010000000000011110, // Bgti (Reg 2) (Imm5 9) (LabelI "then.722.741")
32'b00010000010000100000000000110000, // Addi (Reg 2) (Reg 2) (Imm 48)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000010100000000000000, // J (LabelI "min_caml_print_char")
32'b00101000011000100000000000001010, // Divi (Reg 3) (Reg 2) (Imm 10)
32'b01100100011111010000000000000001, // Sw (Reg 3) (Reg 29) (Imm 1)
32'b01100100010111010000000000000010, // Sw (Reg 2) (Reg 29) (Imm 2)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000011, // Addi (Reg 29) (Reg 29) (Imm 3)
32'b10010000000000000110010000000000, // Jal (LabelI "print_int_sub.328")
32'b00010011101111011111111111111101, // Addi (Reg 29) (Reg 29) (Imm (-3))
32'b01011000011111010000000000000001, // Lwr (Reg 3) (Reg 29) (Imm 1)
32'b00100000011000111111111111110110, // Multi (Reg 3) (Reg 3) (Imm (-10))
32'b01011000010111010000000000000010, // Lwr (Reg 2) (Reg 29) (Imm 2)
32'b00010000010000100000000000110000, // Addi (Reg 2) (Reg 2) (Imm 48)
32'b00001100010000100001100000000000, // Add (Reg 2) (Reg 2) (Reg 3)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000010100000000000000, // J (LabelI "min_caml_print_char")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11111100010111110000000000111000, // Bgti (Reg 2) (Imm5 (-1)) (LabelI "then.728.742")
32'b01001100011000000000010110100000, // Li (Reg 3) (Imm 45)
32'b01100100010111010000000000000001, // Sw (Reg 2) (Reg 29) (Imm 1)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000010100000000000000, // Jal (LabelI "min_caml_print_char")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b01011000010111010000000000000001, // Lwr (Reg 2) (Reg 29) (Imm 1)
32'b00001000010000100000000000000000, // Neg (Reg 2) (Reg 2)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000000110010000000000, // J (LabelI "print_int_sub.328")
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001000000000000110010000000000, // J (LabelI "print_int_sub.328")
32'b01100111111111010000000000000000, // Sw (Reg 31) (Reg 29) (Imm 0)
32'b11111000010000100000000001001110, // Blti (Reg 2) (Imm5 2) (LabelI "then.734.744")
32'b00010000011000101111111111111111, // Addi (Reg 3) (Reg 2) (Imm (-1))
32'b01100100010111010000000000000001, // Sw (Reg 2) (Reg 29) (Imm 1)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b00010011101111010000000000000010, // Addi (Reg 29) (Reg 29) (Imm 2)
32'b10010000000000001110100000000000, // Jal (LabelI "fib.707")
32'b00010011101111011111111111111110, // Addi (Reg 29) (Reg 29) (Imm (-2))
32'b00000100011000100000000000000000, // Move (Reg 3) (Reg 2)
32'b01011000010111010000000000000001, // Lwr (Reg 2) (Reg 29) (Imm 1)
32'b00010000010000101111111111111110, // Addi (Reg 2) (Reg 2) (Imm (-2))
32'b01100100011111010000000000000010, // Sw (Reg 3) (Reg 29) (Imm 2)
32'b00010011101111010000000000000011, // Addi (Reg 29) (Reg 29) (Imm 3)
32'b10010000000000001110100000000000, // Jal (LabelI "fib.707")
32'b00010011101111011111111111111101, // Addi (Reg 29) (Reg 29) (Imm (-3))
32'b01011000011111010000000000000010, // Lwr (Reg 3) (Reg 29) (Imm 2)
32'b00001100011000100001100000000000, // Add (Reg 3) (Reg 2) (Reg 3)
32'b00000100010000110000000000000000, // Move (Reg 2) (Reg 3)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01011011111111010000000000000000, // Lwr (Reg 31) (Reg 29) (Imm 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b10100000010000000000000000000000, // PrintC (Reg 2)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b10100100010000000000000000000000, // ReadI (Reg 2)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b10101000000000000000000000000000, // ReadF (FReg 0)
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b00000100110000100000000000000000, // Move (Reg 6) (Reg 2)
32'b01001100101000000000000000000000, // Li (Reg 5) (Imm 0)
32'b01110000011001010000000001011010, // Bne (Reg 3) (Reg 5) (LabelI "min_caml_init_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100100100001100000000000000000, // Sw (Reg 4) (Reg 6) (Imm 0)
32'b00010000011000111111111111111111, // Addi (Reg 3) (Reg 3) (Imm (-1))
32'b00010000110001100000000000000001, // Addi (Reg 6) (Reg 6) (Imm 1)
32'b10001000000000010110000000000000, // J (LabelI "min_caml_init_array_loop")
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b00000100010111000000000000000000, // Move (Reg 2) (Reg 28)
32'b01001100110000000000000000000000, // Li (Reg 6) (Imm 0)
32'b01110000100001100000000001100011, // Bne (Reg 4) (Reg 6) (LabelI "min_caml_create_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01100100011111000000000000000000, // Sw (Reg 3) (Reg 28) (Imm 0)
32'b00010000100001001111111111111111, // Addi (Reg 4) (Reg 4) (Imm (-1))
32'b00010011100111000000000000000001, // Addi (Reg 28) (Reg 28) (Imm 1)
32'b10001000000000011000010000000000, // J (LabelI "min_caml_create_array_loop")
32'b00000100110000100000000000000000, // Move (Reg 6) (Reg 2)
32'b01001100101000000000000000000000, // Li (Reg 5) (Imm 0)
32'b01110000011001010000000001101011, // Bne (Reg 3) (Reg 5) (LabelI "min_caml_init_float_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01101000000001100000000000000000, // Ss (FReg 0) (Reg 6) (Imm 0)
32'b00010000011000111111111111111111, // Addi (Reg 3) (Reg 3) (Imm (-1))
32'b00010000110001100000000000000001, // Addi (Reg 6) (Reg 6) (Imm 1)
32'b10001000000000011010010000000000, // J (LabelI "min_caml_init_float_array_loop")
32'b00000100100000100000000000000000, // Move (Reg 4) (Reg 2)
32'b00000100010111000000000000000000, // Move (Reg 2) (Reg 28)
32'b01001100110000000000000000000000, // Li (Reg 6) (Imm 0)
32'b01110000100001100000000001110100, // Bne (Reg 4) (Reg 6) (LabelI "min_caml_create_float_array_cont")
32'b10001111111000000000000000000000, // Jr (Reg 31)
32'b01101000000111000000000000000000, // Ss (FReg 0) (Reg 28) (Imm 0)
32'b00010000100001001111111111111111, // Addi (Reg 4) (Reg 4) (Imm (-1))
32'b00010011100111000000000000000001, // Addi (Reg 28) (Reg 28) (Imm 1)
32'b10001000000000011100100000000000, // J (LabelI "min_caml_create_float_array_loop")
32'b00000000000000000000000000000000, // Sqrt (FReg 0) (FReg 0)
32'b10001111111000000000000000000000 // Jr (Reg 31)
};
logic[9:0] in;
integer inst_itr;
integer byte_itr;
integer bit_itr;

initial begin
	CLK = 0;
	inst_itr = 0;
	byte_itr = 0;
	INITIALIZE <= 1;
	@(posedge CLK);
	INITIALIZE <= 0;
	repeat(INST_LEN) begin
		byte_itr = 0;
		repeat(4) begin
			unique case (byte_itr)
				0: in = {1'b1,data[inst_itr][31:24],1'b0};
				1: in = {1'b1,data[inst_itr][23:16],1'b0};
				2: in = {1'b1,data[inst_itr][15:8],1'b0};
				3: in = {1'b1,data[inst_itr][7:0],1'b0};
			endcase
			bit_itr = 0;
			repeat(10) begin
				UART_RX = in[bit_itr];
				repeat(T) @(posedge CLK);
				bit_itr = bit_itr + 1;
			end
			byte_itr = byte_itr + 1;
		end
		inst_itr = inst_itr + 1;
	end
	repeat(100) @(posedge CLK);
	START_EXEC = 1;
	repeat(2) @(posedge CLK);
	START_EXEC = 0;
end

always begin
	#33.3ns CLK=~CLK;
end

endmodule